module main

import code
import ezlang

fn main() {
	code.run()
	ezlang.run()
}


