module ezlang

pub fn run() {
	test_ezlang()
}



