module ezlang

const ezlang_test_path = "./ezlang/test"
