module code

pub fn run() {
	set_edit()
}

