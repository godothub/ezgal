module main

import code

fn main() {
	code.run()
}


